-327
