-3
200
-94
98
167
-97
244
-101
-107
235
-70
-149
-7
136
235
-238
-188
166
-180
50
285
-101
-291
154
-245
-269
51
-164
-127
-145
-83
289
168
65
-42
273
16
91
235
102
-187
-64
-29
187
-228
-239
-272
154
175
99
233
-262
-167
271
-32
179
-296
-144
-39
201
176
220
-121
262
-257
-206
-42
111
-141
80
-202
-17
-234
77
136
-240
-189
256
132
70
-19
-33
-211
-273
-103
274
-84
-169
54
86
-29
3
219
216
-142
271
36
-147
-117
62
-287
-150
-2
-70
-86
105
292
142
216
100
27
-2
-109
-79
288
4
294
-244
298
-262
-43
189
-281
-96
-28
147
-244
-232
-23
235
-265
153
-285
-283
109
-282
286
0
-39
139
160
259
229
184
-176
2
240
109
265
225
74
-235
-166
-98
240
203
263
-111
19
14
-143
101
268
-279
-51
-124
-87
-78
115
95
53
-118
140
-32
-146
-216
222
-196
277
290
-109
-290
-16
-152
-50
110
-217
123
-209
-1
217
86
-86
-137
-87
104
-300
262
87
294
-133
-207
115
-244
-22
149
140
-61
248
81
167
-30
-192
269
165
-16
-187
181
4
27
89
-259
113
155
113
-145
-62
-86
-208
113
-52
40
-164
90
-237
-105
129
32
259
-182
-137
-167
77
190
-36
169
168
42
161
-230
152
176
117
173
-20
-21
-159
141
154
-5
125
-176
-81
63
144
-129
177
88
80
-67
272
233
104
93
81
72
54
140
180
59
-196
-57
-157
-104
-138
239
-48
288
192
-10
-35
282
190
-79
-293
-9
152
217
-279
-203
51
-264
-33
-12
-115
-135
-183
-231
-181
-251
-252
-143
164
254
255
-66
-152
-154
-209
179
62
267
-20
-190
75
86
-39
-41
232
-184
-210
-97
162
276
298
9
140
-103
-172
-187
-266
-139
186
-280
-146
-153
274
-36
77
-293
-9
153
-15
273
-230
-167
-173
-300
226
8
212
-287
-119
180
249
244
32
176
38
141
-108
278
-59
32
-297
-191
-284
-270
-297
-93
156
-212
236
37
-57
212
62
241
-210
-256
-254
268
96
111
-100
266
185
140
279
-212
-9
24
196
130
48
255
-291
-81
217
-146
210
149
-215
240
-41
165
-233
-177
276
-56
188
-115
16
109
-116
219
-133
104
41
-277
-72
-197
-292
-176
92
-134
251
-181
-152
15
-208
-115
57
44
-251
136
-231
-123
173
256
-273
-274
-221
42
-29
-55
123
67
264
177
126
-153
245
289
36
-288
234
-14
222
285
-158
42
187
-167
-11
-163
122
115
9
191
112
297
157
-52
-274
175
-41
254
-260
-82
-292
-286
220
-77
-119
-130
-275
-4
127
-47
293
-143
134
135
-82
269
-251
-99
-218
-130
-193
170
-40
99
-243
-27
274
79
-281
11
48
130
33
51
112
-112
172
-282
49
255
257
69
209
-191
204
63
-238
65
-119
118
164
158
252
-9
-82
-209
-123
172
-259
273
124
227
296
181
282
-245
-155
-153
-238
-235
-245
-127
112
-179
-118
21
-245
-212
-235
-24
-7
-69
52
-141
167
269
-288
80
-142
-38
-215
-73
-126
100
113
-185
-175
-42
291
-170
119
-264
-160
-194
93
252
-50
102
189
-202
118
201
-53
152
-81
186
-131
107
-282
-34
-37
-53
-120
-96
-269
266
-241
251
-59
154
-256
-18
-262
134
117
19
-112
-17
99
-86
221
178
-219
23
81
-184
59
150
286
-213
77
-185
57
94
-102
-137
-107
264
-227
-111
-46
-215
174
247
195
-188
-104
148
-299
-291
-187
-85
20
-187
-170
-173
150
30
64
-118
-72
18
-250
105
51
-208
-230
11
198
40
236
-236
153
161
-79
221
219
38
-203
11
209
-285
74
-256
-110
233
164
125
280
286
-25
-275
-78
-68
-160
-131
-113
246
113
-64
231
48
184
62
-260
47
245
83
271
191
21
-67
19
250
-14
69
1
201
120
-148
-163
109
136
-270
143
-150
-215
-265
87
69
252
51
-178
-204
206
-291
-46
203
-205
-56
-119
-1
51
-120
136
174
245
149
-181
313
-193
222
111
777
686
444
222
777
618
313
-15
75
109
-123
239
-238
-276
116
228
275
196
-128
-166
291
70
-76
217
-33
142
-26
31
218
-227
290
-52
2
217
-139
119
164
-243
192
230
-263
253
-145
-212
87
-280
-15
253
148
-159
-41
-22
34
257
-62
-278
-88
152
152
259
-259
364