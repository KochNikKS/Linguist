-193
222
111
777
686
444
222
777
606
618
364