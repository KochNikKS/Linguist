-327
-936
903
124
829
464
765
-863
163
585
903
200
364
-449
193
200
124
464
765
222
767
767
222
464
606
464
111
777
765
765
765
-200
645
252
124
464
765
111
333
464
333
364
-936
903
124
449
765
449
645
432
200
645
163
585
193
829
422
464
765
-432
464
709
-936
903
124
829
709
-863
163
585
903
200
709
343
829
163
547
124
432
200
903
709
-308
645
585
400
936
645
903
200
765
222
767
767
767
765
-308
-124
709
-449
645
432
709
-124
585
400
308
645
903
618
686
308
449
695
364
-252
163
449
124
464
765
200
829
193
645
585
645
585
400
364
-449
645
829
124
432
200
645
163
585
464
765
-308
124
695
200
765
200
163
765
829
645
400
618
200
364
-903
124
308
124
432
200
645
163
585
464
765
-695
829
163
252
765
200
618
124
765
695
645
829
903
200
765
200
163
765
200
618
124
765
308
193
903
200
364
-193
252
163
936
585
200
765
163
695
765
124
106
343
829
124
903
903
645
163
585
903
464
765
767
364
-193
252
163
936
585
200
765
163
695
765
432
163
829
829
124
432
200
765
193
585
903
643
124
829
903
464
765
767
765
935
767
149
899
364
-193
252
163
936
585
200
765
163
695
765
252
645
903
200
193
863
124
903
464
765
767
765
935
767
149
899
364
319
124
585
449
920
364
-936
903
124
829
464
765
-863
163
585
903
200
364
-449
193
200
124
464
765
222
767
767
222
464
606
464
111
777
765
765
765
-200
645
252
124
464
765
111
333
464
777
364
-936
903
124
449
765
449
645
432
200
645
163
585
193
829
422
464
765
-432
464
709
-936
903
124
829
709
-863
163
585
903
200
709
343
829
163
547
124
432
200
903
709
-308
645
585
400
936
645
903
200
765
222
767
767
767
765
-308
-124
709
-449
645
432
709
-124
585
400
308
645
903
618
686
308
449
695
364
-252
163
449
124
464
765
200
829
193
645
585
645
585
400
364
-449
645
829
124
432
200
645
163
585
464
765
-308
124
695
200
765
200
163
765
829
645
400
618
200
364
-903
124
308
124
432
200
645
163
585
464
765
-695
829
163
252
765
200
618
124
765
695
645
829
903
200
765
200
163
765
200
618
124
765
308
193
903
200
364
-193
252
163
936
585
200
765
163
695
765
124
106
343
829
124
903
903
645
163
585
903
464
765
767
364
-193
252
163
936
585
200
765
163
695
765
432
163
829
829
124
432
200
765
193
585
903
643
124
829
903
464
765
767
765
935
767
149
899
364
-193
252
163
936
585
200
765
163
695
765
252
645
903
200
193
863
124
903
464
765
767
765
935
767
149
899
364
319
124
585
449
920
364
